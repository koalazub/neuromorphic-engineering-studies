module  HelloWorld;

initial
  $display("oi oi");

endmodule
